																																																																																																																																																																																																																																																														****************    ****																																																																																																										****************																																																																																																																																																																																																																																			      																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																				  																																																																																																																																																																																																																																																																																																																																																																																																																																																			   																					































































































































































































																																																																																														









																																																																																																																																																																				  							  

                    																																											          																																																																																																																																																																																																											  					

















































   















































   																																																																																																																																																																																											























																																																														   																																																																																																																																																																																																																																																																																																																																																																																																																																																																																				







   








 
  																																																																																																																																																																																																																								







        















    



        																																																																																																																																																																																																									  																		



 



          


 


              																																																																																																																																																																				                            																																																																																																																																																																																																																																																																																																																																																																																																	

























































































































 

 

 

 














































































































































































































																																																																																																																																							    																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																										
   
																																																																						  













																																																																																																																																																																																																																																																								





  





  






 






 																																																																																																																																																																																																																																																																																																																																																																																				     							


									     		  																																																																																											





																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																								































																																									   																															


																																													  																																																																																		
   

    																																																						**********************  ******* *******         ******* ******* ****************                                                                                                                                                                                                        ******  *****           ******  ******  *****         																																																																																																																                                                                                                                                   ..      ....      ....      ....      ....      ....      ......    ....      ....      ....      ....      ....      ..                ..................  ..........................................................................................................................................................................................................................                                                                                                                    .............................................................................................                                                                    .......................................................................................................................                                                                                                                                                                                                                                                                                 ...................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................    .............................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                      ...............................................................................................................................................................................................................................................................................................................................................................................................................................               .........................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ......................................................................................................................                                                 .................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             