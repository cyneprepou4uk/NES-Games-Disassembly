                                                                















                                																																																																																																																																																																																																																																																																																			      																															      																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																								



																																																																																																																																																																																																							   																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																					     																																																																																																																																																																																																																												





																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																										*********************************************************************************************************************************************************************************************************************************************************************************************************************************************











                                   																																																																																																																																																																																																																																																									      																																																																																						































































































































































																																																																																																																																																																																																																																																																																																																																																																				        																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																			             																																																																																																																																																																																																																																																											













 
























































    



																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																										                      ..  ..      ..........            ..                                                          ...............................................................................................................................................................                               .................................................................................................................................................................................................................................................................................................................................................................................................                                                                                                                                           ............................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      