J               																																																																																																																																																																																																																																																								******************																																																																																																																																											








			******************																																																																																																												 																																																																																																																																																																																																																																																																																																																																																																																      																																										  	                       																																																																  																																																																																																																																												

********************************																																																																																																																	                													  																																																																									

																																						  																					           																																												

																																																																																																																																																											********																										                        													  																																																																																																																									       																						  																																																																																																																																																																								 																																																																																																																																																																									            

									            																			******************************************                    ***********************************************************************************************                           ****************************************************************          *******************************************************************************        *********************************************************     *****    *******                 *********************************













  





























********************************************************************************************************               ***************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************** ************************************************************************************************************************************																																																																																																								



																																																																																																																																																																																																																																																																																																																																					   																																																																																																																																																																																																														  







  

  







																																																		 																										******  ******  ******          ******  ******  ******          ******  ******                  										


 


 


                    																					
























            																																																																																						      												             																																																											      					      																																																																																																																																																																																    																																																																																																																												    																																						**************																																																																																																																																																		 





 																																																																															 																																																																																																																																																																																																																																																						**********																																																																																																							****  																																																				                					 








































																																																																																																																																																		





















***********************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************																																																																																																																																																																																																																										   																											 																																																																																														  

 



       







































																																																																																													  																			


																																																																																																											  																																																																																																																																																																																																																																									  																																																																																																																			                          																																																																	



																																																																																																																																		


						 																																																																																																																																																																																																																																																																					


																																																																																																																																																									                .               .               .               .               .               .               .                                                                                                                                                                                                                           ........................                                                                                                                                                                                                                                             ..........  ..........  ..            ........    ..    ......          ........  ..                    ........  ..    ......        ..........                                                                                                               ....................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................     .........................................                 .......................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................           ............................                        ..........                                                                                                                                                                                                                                                                                                    ....  ......  ................  ......................    ..      ....    ......  ..    ..                                                                                                                         