



























































********************************************************************































































 

































































 










  












 










  





















     












































    











																																																																																																																					   																																																																																																																																																																																																																							  																																																																																																															               																																																																																																																																																																																															                           																																																																																																																																		    																								    																																																																																																																																																																																																																																																																																																																													           																																																																				                                                    																																																																																																																										                                                                                							                                                                     																																																																																																																																																																																																																																																																																										   																							    																																																																																																																																																																																																																																																											                        																																																																		     																																																																																																																																																																																																																																																																																																																																																																																																																																																																																								   																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																          																																																																																																																																																																																																							*******************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************               *****************************         ****************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************  


 


 


 






 


 


 



























































































 

 



















































																																																																																																																																																																																																		   																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																								      																																																																																																																															      ......................................................................................................................................................................................................................................................................................                                                                   .............................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................  ...........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                                                        .....................................................................................................................................................................................................................................................................            ......................................................................................................................................................                                                                                                                                                                                                                                                                                                                                  